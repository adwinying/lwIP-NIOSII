��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O����w��=�3�n����0:��q�q��%�J�`���l�d6��p�y~ �z8`���K�<��"�em²�݌�x@0�^ W�wK�߿�=��:1�ʅ���*h�1g�^O�v��z�sYt�}��Δ��!���@ݻ]0��1�d�Tz:=܉
��-���9��`=_�x&�/H��[(���d=����`�X���}U*^Z7~Q�U����jp��;����T
-���hU��cͧ\b,ܕ�*��l�O{i{��hE̿���J� �l��X��)�t��#�1����\Q���^	r]���ͣ@,�ea%0ʨ$m�
kg�(a3_�4w���Ź�0?�*�я&��h�-� � F(��p�c������u��t�L��EmdH}��JUʥ�'��`�ni��+�vu>.�<��[v�W�M��'�UH,���]�4�mѻ�n�DXG9u�ST@/�8�$�Ch7��gW)�6P�<#XǮ9Z�#X�o�1A����������o�E̩�mB�1�_xc�+ �Q��s����;���{R�[�Xد��h���ku?8������%{jLu�:����2OcO�����_{$=?�}�g3�o(d\��|��-�i6�]6)�V�DN��kǕ�Av�;<{�e�`�@�g��q)�~gc�׽�I������Y��uVG�Ĳ����8������>o�Em���.۝��/y�X4f�Η;��;�E�̃nh��_�bug����֠����xL�v�rnK�������f8�i��43\��o��Wd��*&�B��X
}�O��I�c�1S�l�̬�Y��C�d��}��^�y�U�B��G��$,?�YݕDSM��i&�]{�jE�g�j�!OW�W����'�o	�J�dԨ�0Wm$4��9��n�4C�ҍA����m�H�\�P�����p�H�:}��x���܎(n���O5�
q���ٓV\&�����{E$EKr>t<xa�Dj	B�o�Ќ�:����g�d1����Dl�J��r����B�����8�>ᝄ����rN�r���a���{=4���1�z���xr�%�K�"{��e#v��ڜm�Q9,ugs�ɢ�{�$�)��}8#�	8";i�!�ɓ1Wh���(����a��}[��f1��������Ψ!gFCk��mnE�^18YE5�b�tg
��i��{.b2�1#m�]l���$�D(q����]'1ws�17��O��2�(��W*�k�@��ӂF�|8�Q:��K@5��`A�,0f�����>,iw�Z���-pUǇI��t��OP7�D��������o"i]���U^E#��&��jK<���YU7&M��_��JG�(%$q��m�r�����n{W�wLk&���v�EC*#�p�2 �Ӆ>u8�~?أ�K���"���*�53����=��Tq�ł8KV_{��J����7�ЪU��@�y��OEu�8@��>9������N�*�F�R��T&!X �CݼLV����?�MH5���\�"�S��Ak�)�Zr�
��(��6@Y�-!�Y�d�����n��>��5�`��#��5������e�/_\��X���t�R���#�-#B��,��}�k \�o:#��� �'��+0���"�OF�-���]�\�gz|k�T�ՠ�˭nl_ x�'��}���Zi=e�8�����u98O=SЅ���4��nE���ΆD9�Ig�Z7��k���92�����ੇE�4^�b`�Ocζ�)�����y#a�} M_���a�r�z�yI�[*�{�<L�F1J�m�=%����r��,ehڗ�R��iC���3s�ѿ^� �����{�s��Ɓ*�M�yP������?EIŽ%� Ӄ*D[�.�}>7=6���9S�B��Y'��;�~p��J݆v�O�sp5�Ф��:�[蒱!w0�A�A쀟���W|&*@��:Yg-S�.�0�	 �Z�#A��\:VJ4�ak9��<zBV�����`�k���%Zf�AWh��b<���gm`�f/Y�l�7T!���.޸�4�z\��0��������&e)���?��/ܴ�ƒT$1�nm�w�0Z:���8����4h�y�x�䥝�ה�D�$������sw�S�,
R�m�"���(в�����Ԥ$ќ]���J���y�˕^�a�$ZH���3\I:DR���ʓ>y������,=�e��~��=��^��B�v�8s�5�=�e#�g�3��F;���v��}�O۵5�<!�|�S� 3���_ؚ�{*�]��v�̄�A�)�땲C �����*	�7.ɘ��X��h����{}���b���4�HF@I����+�R:�陵������N�'^���UCw����~"�����PbB-�@�5?���� �P�=����E5)m�99�B3S}*��d6�`0^�?�!>� �^5�j7� CݴOť&B �b ֫�r�ˤ�P��l��$/�c����<�*�t�O��O�O�(=��m��?��EqR!X�T�u��f���ٵ��B,Ɗ����%8_c�<H�0ƕ��_����������s4I�(�G�(ˡ2rl1���1�PO�Kw�O����B�����.����c|�<m��]JNS#�2�� ����Lu�nP���\u|��r�)�\W}�	頻 ���8�A/6WK������K(�8S�_���%�A��u
Vǋ�R�]I��<\_���Mf��1��+/��B��k-��ev)���]�^'��)�����9c�a�e�����kO�D�7I��FE �%��_e���ٴv�9&Ŷ��HW�L]�<��Ѕ�u�M� ���H��=��ي�%_P�&�c�е�|3zr�p�����QS�&#���,t��ɓ�{��˙[��j�.j�֬�1�/~:���2�Nb/��߱�0{���lʐ�$B �V(�\�ulNysftY��k���8X��c�t�;f�+݉���%��t�� f����q�Y���!���] ��-��8{*�� \u� M�ҋoPxYVk��EWU��KuŦ�b�(�fԇ���7�R.�5��oMl�	�C&�+>	�2W�x�E
ϱ��m�ѕ+GT�QO��|o.�C������LG"1o�24����/*E�z^�/��%��~����HpV�5���
.	��D�i'RC.P	��6V[�),�{I�w�����v��z"���/�I��ʜ��%F#�C>�m�7U��f�K�@�Z�a��r�11���*�������_�=y*m���}�uǳ�|Hl0�Vt,������U�4���F��0d������IB�����:;u�?^XoDɁ��r��.�����.D���`�h0��(Iܒ����϶+�-��L�K J�d��7v�t�tJ�e�K��+��6�u��ټDN����V��q�g�o&����=�_W?�0�V��e��3�$��Q-̘no1�� � #	ָ޾�����О���$[ssRZ��T'�]�?2`�ޚ�ڋ^|�d�p�>2��S��wUy�"i�� U���L6Z36���#���5i��M����r�$�Eոe�UG���>����)�h��Yh�|j�L�H9����yE�O�$܉WJ<��Ժ����u����̺P*�	��"�3u`�ՠ�_�DL�#���S(D�f*\C�
�������>5�IMU�!y ��^������	G{��C3�6���n�'	6�/\JCC��S�~M��L!Xk-����Ԃx�҂.^HrT1U������^���!^d�c��J@`[}�����sZ�tT>�P6<-ҫmnK����ڳ0�m��h1��t��tL\��%b�6w�a��wtM�q����j��l�'J-*9BV�0�H���FE�AB���3ts���"ֹʱJklQ��5#�Ϻs�Y�V�m�	'ܶLg���X0{��k_9��ǎ���3��M
�݄h�)��u �6�JBR�. !淫��Csu����їg&�=�_b�gu��Q��{����dץ����{�<���d|d��d=jK�4b"{�.&�?�w���k�\�q?�X�y����c�����R�~�XǊ��P!xp^N�z}.	�כ��"М�Q�5n&���]���n�K�^D�mz{��)f��]���]�p%s�7��E�UM�,�(�̻K�=뺡8�ْæ��
f�-���۾��^�R)QV��ո.�Qx��&!��>�K����tÚ�>������|���4O�?`�N{`�g���v���_캁���6ucd��d*��� �-Vo��1Ӎ�8Ъ#Ԅm;N��	Q'{Ӝ�Ň;g{�b���Y0�ڨ��w������<ߛ�g��|�]ٌє�\���@�|��(��4��ZrV�Ehnůk���O�a�TL��W�[�M�d!o�(�<0SkB���X��/C�z�N����H�5��Ky�����~�伣��;y�C9��{~Ư+�Z.&��t��n��v�O_x�~�A�ߨ��I54.��W!��A
��*Z��"��![����\�ݱ')#$6��o�5ҰB̭���6�Us���A;�X'{�oA�Gm�\j�p���wd�5���Jr���l�a��$�DW�q���Z�`����l�}j�O��~���j��,�e�j� �j�f�͔\]5X]�'�&��7�1��X^-d�񷌖�An�9	��>����HtV���0�� {El�_�)Vow�����.P}'����o�;�Ա���l�z6R:���m5g�ɤyb���|��G���&1��6��0��+���X�;'�e=��irqgѨ���U�%���o.g����� �tz.5�j[U�����3����@ �������r!�F�S#q��Wuϥ��{�4s��	�8���G���;����ʫx�<��&vmeL��S���V�;$��9T@�Ǟm'5�V"V������K$���N�e��������쐢]���؅4_���5��0҂��x!�m�� )]v�A���Pe�DD9S�D��l�/�C��,�fcG�c,X�QvZ	���&J!��pyH�.Nr�3J�1z�)�eR�L3��k��l���~A��a�7\?�➨&����	�M ��̩����@�;soAI�6�SYv�߸a_*~7��a
{i��(�.�H"��\"��r�kk�pXM����U��g15g@�g��	��k��ݗ�{��dm%@��3��
�'lw�hpzYl���Y�/��"û�n��1<�3�Q!��e�1�P��] �I�.��n�|�z���h�DdR�s���?��lix���K�6b��c���Si���S��!��ސ���·�e3����f��ڋ�ڡ�.��;w*����U��O�B�n�:������̈,*`�G�ޘ�2��¡�z۪�-cIS%�yn�V�����nCH%=4��{������A]��̤	�/�;��]z�ʿ���o��]���AOI=	��e]��G�NVӥ��G�@��n�}yM1.��)]z����o%���'�`���<[�ť��;e|�w����# ���Y86��y����:���K\i�wb��&�_�<�|���N�AWr��֧qr>w_��� ���Ht����ٸ{~x�3�E��_Yo �@ږ5�7�/���JV��������҂���h����^�'ܵ��$㨒�S �R@�A*�H6��ǖL��R�_u��h����1�2�"��1���+u&���) �ҵ��>�#V]���+�kpu5I�J(ЎL:��|[�6�_䉳�_$el�p����WbF�(�M
�΃�/�RDX���^�0H�_8n�/�l4p�4��@���a���j���1B��̪d��_=��������t�NdP�ǅ��%gdj[,���ch6yI�4?��%=.Z��قxWr�ߤ�b�-�@����
�;��p�̿ŕ7�%*`Z�rK~F�&]�&j�k��Y�BX�3�hcp¸VtZ� ���>P��G)�� Ф��{9��p�PlY¡�Nn�o�rV�2�%�S��%�S�ҧ=�E0Y�p(yP�����]�~I;K�����Q���oX�k8���������i<���r9��n&v�P�լ��͜�˂���+�='��-���